
library IEEE;
use IEEE.std_logic_1164.all;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY REGFILE IS
PORT(
	RD1: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    RD2: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    WR1: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    DATA: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    W_SEL: IN STD_LOGIC;
    CLK3: IN STD_LOGIC;
    OUT1: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    OUT2: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END ENTITY;

    
ARCHITECTURE BEH OF REGFILE IS
TYPE MEM IS ARRAY(15 DOWNTO 0) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL MEMORY : MEM:=(
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000010",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000");


BEGIN
PROCESS(clk3)
BEGIN
if (rising_edge(clk3)) then
	IF(W_sEL='1') THEN 
     	MEMORY(CONV_INTEGER(WR1))<=DATA;
    else
        OUT1<=MEMORY(CONV_INTEGER(RD1));
    	OUT2<=MEMORY(CONV_INTEGER(RD2));	
    END IF;
end if;
END PROCESS;
END BEH;